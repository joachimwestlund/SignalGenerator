* AD8021 Spice Model             
* Description: Amplifier
* Generic Desc: 250MHz very low noise op amp
* Developed by: TRW
* Revision History: 08/10/2012 - Updated to new header style
* 4.0 (10/2001)
* Copyright 2001, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.
* Use of this model indicates your acceptance with the terms and provisions in the License Statement
*
* BEGIN Notes:
*
* Not Modeled:
*       distortion is not characterized       
*       disable is not characterized
*
* Parameters modeled include:
*       open loop gain and phase vs. frequency
*       output voltage 
*       Common Mode Rejection
*       input common mode voltage range
*       slew rate
*	Voltage noise
*	Current noise
*	Output current to supplies
*
* END Notes
*
* Node assignments
*                   non-inverting input
*                   |    inverting input
*                   |    |    positive supply
*                   |    |    |    negative supply
*                   |    |    |    |    output
*                   |    |    |    |    |     Ccomp
*                   |    |    |    |    |     | 
.subckt AD8021      1    2    99   50   45    10

***** Input stage

Rc1 99 4 rmod 1190
Rc2 99 5 rmod 1190
Q1 4 1 6 nbjt
Q2 5 3 7 nbjt
Re1 6 8  rmod 1128
Re2 7 8  rmod 1128

Ibias 8 50 840u

***** Input Error Sources

eos 2 3 poly(2) 30 98 64 98 39.6e-3 1 1e-3
gnoise1 98 1 33 98 1e-4 
gnoise2 98 2 33 98 1e-4

Cin+ 1 0 2pF
Cin- 2 0 2pF
Rin 1 2 10Meg

****** CMR Stage

Gcmrr 98 64 97 98 13n
Rcmrr 64 65 rmod 1e6
Lcmrr 65 98 1.59

****** Gain Stage & Dominant Pole

Rgain1a 98 10 rmod 1.3263Meg
Ggain 98 10 4 5 13.48m
Cgain1a 98 10 2e-12

Dpvc 10 80 diode
Vpvc 99 80 2.28

Dnvc 81 10 diode
Vnvc 81 50 2.68

****** Second Pole

Ggain2a 98 13 98 10 0.01
Rgain2a 98 13 100
Cgain2a 98 13 0.80p


****** Reference Stage

Eref1 98 0 poly(2) 99 0 50 0 0 0.5 0.5

Eref2 97 0 poly(2) 1 0 2 0 0 0.5 0.5

****** Voltage noise stage

rnoise1 39 98 7.3e-4

vnoise1 39 98 0
vnoise2 31 98 0.75
dnoise1 31 39 dn
fnoise1 30 98 vnoise1 1
rnoise2 30 98 1

****** Current noise stage

rnoise3 32 98 0.166e-3
vnoise3 32 98 0
vnoise4 34 98 0.545
dnoise2 34 32 dn
fnoise2 33 98 vnoise3 1
rnoise4 33 98 1

****** Output Stage

Dout1 13 11 diode
Dout2 12 13 diode
V1 11 44 -0.884
V2 44 12 -0.884

Vo1 91 99 0
Go1 91 44 13 99 15.823
Go2 44 51 50 13 15.823
Vo2 50 51 0

Rout1 91 44 .0632
Rout2 44 51 .0632

Vout 44 45 0

Fout 98 72 Vout 1
Diout1 72 74 diode
Diout2 73 72 diode
Viout+ 74 98 0
Viout- 73 98 0

Fsy+ 99 0 poly(2) viout+ Vo1 6.25e-3 1 1
Fsy- 0 50 poly(2) viout- vo2 6.243e-3 1 1


.model rmod RES(t_abs=-373)
.model diode D(IS=1e-15)
.model nbjt npn(bf=56)
.model dn d(kf=1e-13,af=0.55)
.ends
                      





